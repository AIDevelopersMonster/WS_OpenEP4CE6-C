// ------------------------------------------------------------
//  Module     : fmq
//  Project    : Buzzer Signal Generation
//  Description: 
//    Модуль генерирует выходной сигнал для управления 
//    пищалкой (buzzer). Сигнал меняется с определенной частотой.
//    Для работы требуется тактовый сигнал (clk) и активный сигнал 
//    сброса (reset). Сигнал на выходе меняет свое состояние через
//    каждые определенное количество тактов (по счетчику).
//
// ------------------------------------------------------------

module fmq(
				clk,        // Тактовый сигнал
				reset,      // Сигнал сброса
				out         // Выходной сигнал
           );

input clk;               // Входной тактовый сигнал
input reset;             // Входной сигнал сброса
output out;              // Выходной сигнал, который будет управлять пищалкой

// Регистр для отсчета тактов
reg [23:0] cnt;           // 24-битный регистр счетчика

// Счётчик увеличивается с каждым тактом и сбрасывается, когда достигает значения 24'hFFF
always @(posedge clk or negedge reset) begin
    if (!reset)               // Если сигнал сброса активен, счетчик обнуляется
        cnt <= 24'd0;
    else if (cnt == 24'hFFF)  // Если счетчик достиг значения 24'hFFF
        cnt <= 24'd0;         // Сбрасываем его
    else
        cnt <= cnt + 1'b1;    // Иначе увеличиваем на 1
end

// Регистр для выхода
reg out_reg;

// Переключаем выходной сигнал на основе счетчика
always @(posedge clk or negedge reset) begin
    if (!reset)              // Если сигнал сброса активен, выходной сигнал устанавливается в 1
        out_reg <= 1'b1;
    else if (cnt == 24'hFFF)  // Когда счетчик достигает 24'hFFF, инвертируем выходной сигнал
        out_reg <= ~out_reg;
end

// Присваиваем выходному сигналу значение из регистра
assign out = out_reg;

endmodule

// ------------------------------------------------------------
//  Module     : sel_4
//  Project    : 4-digit multiplexed display driver
//  Description: 
//    Этот модуль управляет 4-значным дисплеем с помощью мультиплексирования. 
//    Он управляет выбором активной цифры и отображает её на 7-сегментном дисплее.
//    Входной сигнал "number" представляет 16-битное число, которое разбивается на 4 цифры,
//    и каждая из этих цифр отображается поочередно на дисплее.
//    Время переключения между цифрами составляет 10 миллисекунд.
// ------------------------------------------------------------

module sel_4(
    input clk,           // Тактовый сигнал
    input nrst,          // Сигнал сброса (активный низкий)
    input [15:0] number, // 16-битное число для отображения
    output reg [3:0] sel,  // Выбор активной цифры
    output [6:0] seg      // Управление сегментами 7-сегментного дисплея
);

    reg [3:0] data;       // Хранит текущую цифру для отображения
    reg [31:0] count1;    // Счётчик для задержки
    reg sel_clk;          // Тактовый сигнал для выбора активной цифры

    // Модуль для задержки 10 мс
    always@(posedge clk, negedge nrst)
    begin
        if(!nrst) begin
            count1 <= 0;
            sel_clk <= 0;
        end
        else if(count1 == 50000) begin  // Задержка 10 мс (при тактовой частоте 5 МГц)
            count1 <= 0;
            sel_clk <= ~sel_clk;  // Переключаем состояние тактового сигнала
        end
        else begin
            count1 <= count1 + 1;  // Увеличиваем счётчик
        end
    end

    // Мультиплексирование цифр
    always@(posedge sel_clk, negedge nrst)
    begin
        if(!nrst) begin
            sel <= 4'b0001;  // Начинаем с первой цифры
        end
        else if(sel == 4'b1000) begin
            sel <= 4'b0001;  // После последней цифры начинаем сначала
        end
        else begin
            sel <= sel << 1;  // Сдвигаем влево, чтобы выбрать следующую цифру
        end
    end

    // Выбор соответствующих 4 бит данных для текущей цифры
    always@(*)
    begin
        case(sel)
            4'b0001: data = number[3:0];   // Первая цифра (младшие 4 бита)
            4'b0010: data = number[7:4];   // Вторая цифра
            4'b0100: data = number[11:8];  // Третья цифра
            4'b1000: data = number[15:12]; // Четвертая цифра
            default: data = 0;             // По умолчанию сбрасываем данные
        endcase
    end

    // Модуль для управления сегментами дисплея
    seg_7 output_seg(
        .data(data),  // Текущая цифра для отображения
        .seg(seg)      // Выходные сигналы для сегментов
    );

endmodule

// ------------------------------------------------------------
//  Module     : seg_7
//  Project    : 7-segment display decoder for 4-bit data input
//  Description: 
//    Этот модуль преобразует 4-битный двоичный вход (data) в управляющие сигналы для
//    7-сегментного дисплея. Каждый входной символ (0-15) отображается на дисплее 
//    соответствующей цифрой или буквой, где 0 - это отображение цифры 0, 1 - цифры 1 и так далее.
//    Сигнал "seg" будет управлять сегментами дисплея, где 0 активирует сегмент, а 1 - деактивирует его.
// ------------------------------------------------------------

module seg_7(
    input [3:0] data,  // 4-битный входной сигнал (данные от 0 до 15)
    output [6:0] seg   // 7-битный выходной сигнал для управления сегментами дисплея
    );
    
    reg [6:0] seg2;  // Временный регистр для хранения данных сегментов

    assign seg = ~seg2;  // Инвертируем значение, так как для активного сегмента на дисплее требуется логический 0
    
    // Преобразование 4-битного входного значения в соответствующие управляющие сигналы для 7-сегментного дисплея
    always@(*) begin
        case(data)
            4'h0: seg2 = 7'b1111110;  // 0
            4'h1: seg2 = 7'b0110000;  // 1
            4'h2: seg2 = 7'b1101101;  // 2
            4'h3: seg2 = 7'b1111001;  // 3
            4'h4: seg2 = 7'b0110011;  // 4
            4'h5: seg2 = 7'b1011011;  // 5
            4'h6: seg2 = 7'b1011111;  // 6
            4'h7: seg2 = 7'b1110000;  // 7
            4'h8: seg2 = 7'b1111111;  // 8
            4'h9: seg2 = 7'b1111011;  // 9
            4'hA: seg2 = 7'b1110111;  // A
            4'hB: seg2 = 7'b0011111;  // b
            4'hC: seg2 = 7'b1001110;  // C
            4'hD: seg2 = 7'b0111101;  // d
            4'hE: seg2 = 7'b1001111;  // E
            4'hF: seg2 = 7'b1000111;  // F
            default: seg2 = 0;  // По умолчанию выключаем все сегменты
        endcase
    end
    
endmodule
/*

Пояснения к коду

Входные и выходные сигналы:

data: 4-битный входной сигнал, который может принимать значения от 0 до 15 (0x0 - 0xF).
 Эти данные будут интерпретированы как цифры или буквы для отображения на 7-сегментном дисплее.

seg: 7-битный выходной сигнал, где каждый бит управляет соответствующим сегментом 7-сегментного дисплея (от A до G). 
Логический 0 включает сегмент, а 1 выключает его.

Инвертирование сигнала:

assign seg = ~seg2;: На дисплее для активных сегментов требуется логический ноль. 
В коде для активного состояния сегмента устанавливается 0, а для неактивного – 1. 
Поэтому перед выводом на дисплей происходит инвертирование сигнала.

Логика отображения цифр:

Внутри блока always@(*) используется конструкция case, которая проверяет значение входа data
 и на основе этого генерирует управляющие сигналы для каждого сегмента дисплея. 
 Например:

Когда data равно 4'h0 (0 в шестнадцатиричной системе), на дисплее будет отображаться цифра 0 (seg2 = 7'b1111110;).

Когда data равно 4'hF (15 в шестнадцатиричной системе), на дисплее будет отображаться буква F (seg2 = 7'b1000111;).

Пояснение конструкции языка:

case: Это конструкция языка Verilog, используемая для выбора одной из нескольких альтернатив 
в зависимости от значения выражения (в данном случае, значения переменной data). 
Это аналог оператора switch в других языках программирования.

assign: Это оператор, который используется для присваивания значений выходным сигналам или регистрам в Verilog. 
В данном случае используется для инвертирования сигнала перед выводом на дисплей.

Инвертирование (~): Оператор инвертирования в Verilog. Он меняет все биты на противоположные. 
Здесь он используется для инвертирования выходного сигнала, чтобы соответствовать логике работы дисплея.

Как использовать этот модуль:

Этот модуль можно использовать в проекте для управления 7-сегментным дисплеем, где вам необходимо отображать
 цифры или буквы на основе 4-битных данных. 
 Например, если вы хотите отобразить число, передавайте его в data, и соответствующие сегменты
 будут управляться автоматически.




*/
/*
 * Модуль: LED_4
 * Описание: Модуль для управления 4 светодиодами (LED) с использованием FPGA.
 * Реализует последовательность переключения светодиодов с использованием делителя тактовой частоты.
 * Светодиоды переключаются поочередно каждые несколько тактов.
 *
 * Входы:
 *  - nrst: сигнал активного низкого сброса (reset).
 *  - clk: основной тактовый сигнал.
 *
 * Выходы:
 *  - led: 4-битный сигнал для управления светодиодами (LED).
 *
 * Автор: Alex Malachevsky
 * Дата: 23.11.2025
 * Версия: 1.0
 */

module LED(
    input nrst,          // Сигнал активного низкого сброса (reset)
    input clk,           // Входной тактовый сигнал (clock)
    output reg [3:0] led // Выходной сигнал для управления светодиодами (LED)
);

    reg [31:0] counter;  // Счетчик для делителя тактовой частоты
    reg clk2;            // Разделенный тактовый сигнал для обновления светодиодов
    reg [7:0] i;         // Счетчик для последовательности светодиодов

    // Логика делителя тактовой частоты: генерирует сигнал clk2 с частотой ниже, чем clk
    always @(posedge clk or negedge nrst) begin
        if (!nrst) begin
            counter <= 32'd0;  // Сбрасываем счетчик при активном низком сбросе
            clk2 <= 0;         // Обнуляем разделенный тактовый сигнал
        end else if (counter == 1250000) begin
            counter <= 32'd0;  // Сбрасываем счетчик, когда он достигает 1250000
            clk2 <= ~clk2;     // Переключаем clk2 на противоположное значение (делаем его периодическим)
        end else begin
            counter <= counter + 1;  // Увеличиваем счетчик при каждом такте
        end
    end

    // Управление светодиодами, обновляемое с помощью сигнала clk2
    always @(posedge clk2 or negedge nrst) begin
        if (!nrst) begin
            led <= 4'd0;  // При сбросе светодиоды обнуляются
            i <= 0;       // Сбрасываем счетчик последовательности
        end else begin
            case (i)  // В зависимости от значения i выводим разные паттерны на светодиоды
                0: begin 
                    led <= 4'b0001;  // Включаем первый светодиод
                    i <= i + 1;      // Переходим к следующему состоянию
                end
                1: begin 
                    led <= 4'b0010;  // Включаем второй светодиод
                    i <= i + 1;      // Переходим к следующему состоянию
                end
                2: begin 
                    led <= 4'b0100;  // Включаем третий светодиод
                    i <= i + 1;      // Переходим к следующему состоянию
                end
                3: begin 
                    led <= 4'b1000;  // Включаем четвертый светодиод
                    i <= 0;          // Возвращаемся к первому состоянию, чтобы цикл повторился
                end
            endcase
        end
    end

endmodule

/*
 * Пояснения:
 * 1. Сигналы и переменные:
 *    - `nrst`: активный низкий сброс, используется для сброса состояния модуля и сброса всех регистров.
 *    - `clk`: основной тактовый сигнал, который используется для обновления состояния системы.
 *    - `led`: 4-битный выходной сигнал для управления 4 светодиодами.
 *    - `counter`: 32-битный счетчик для деления частоты тактового сигнала `clk`.
 *    - `clk2`: разделенный тактовый сигнал, частота которого ниже, чем у основного сигнала `clk`.
 *    - `i`: 8-битный счетчик для индекса текущего состояния последовательности светодиодов.
 *
 * 2. Делитель тактовой частоты:
 *    - С помощью счетчика `counter` генерируется сигнал `clk2` с более низкой частотой.
 *    - Сигнал `clk2` используется для управления обновлением состояния светодиодов.
 *    - Когда счетчик достигает 1250000, сигнал `clk2` переключается, обеспечивая низкочастотный сигнал для управления светодиодами.
 *
 * 3. Управление светодиодами:
 *    - Светодиоды переключаются поочередно. Каждый новый светодиод включается через один цикл `clk2`.
 *    - Когда значение счетчика `i` достигает 3, оно сбрасывается, и цикл повторяется.
 *
 * 4. Принцип работы:
 *    - Когда модуль сбрасывается (`nrst` = 0), все регистры (включая светодиоды) сбрасываются в нулевое состояние.
 *    - После сброса светодиоды начинают поочередно включаться и выключаться с использованием делителя тактовой частоты.
/*
 * Модуль: LED_4
 * Описание: Модуль для управления 4 светодиодами (LED) с использованием FPGA.
 * Реализует последовательность переключения светодиодов с использованием делителя тактовой частоты.
 * Светодиоды переключаются поочередно каждые несколько тактов.
 *
 * Входы:
 *  - nrst: сигнал активного низкого сброса (reset).
 *  - clk: основной тактовый сигнал.
 *
 * Выходы:
 *  - led: 4-битный сигнал для управления светодиодами (LED).
 *
 * Автор: [Ваше имя]
 * Дата: [Дата]
 * Версия: 1.0
 */

module LED_4(
    input nrst,          // Сигнал активного низкого сброса (reset)
    input clk,           // Входной тактовый сигнал (clock)
    output reg [3:0] led // Выходной сигнал для управления светодиодами (LED)
);

    reg [31:0] counter;  // Счетчик для делителя тактовой частоты
    reg clk2;            // Разделенный тактовый сигнал для обновления светодиодов
    reg [7:0] i;         // Счетчик для последовательности светодиодов

    // Логика делителя тактовой частоты: генерирует сигнал clk2 с частотой ниже, чем clk
    always @(posedge clk or negedge nrst) begin
        if (!nrst) begin
            counter <= 32'd0;  // Сбрасываем счетчик при активном низком сбросе
            clk2 <= 0;         // Обнуляем разделенный тактовый сигнал
        end else if (counter == 1250000) begin
            counter <= 32'd0;  // Сбрасываем счетчик, когда он достигает 1250000
            clk2 <= ~clk2;     // Переключаем clk2 на противоположное значение (делаем его периодическим)
        end else begin
            counter <= counter + 1;  // Увеличиваем счетчик при каждом такте
        end
    end

    // Управление светодиодами, обновляемое с помощью сигнала clk2
    always @(posedge clk2 or negedge nrst) begin
        if (!nrst) begin
            led <= 4'd0;  // При сбросе светодиоды обнуляются
            i <= 0;       // Сбрасываем счетчик последовательности
        end else begin
            case (i)  // В зависимости от значения i выводим разные паттерны на светодиоды
                0: begin 
                    led <= 4'b0001;  // Включаем первый светодиод
                    i <= i + 1;      // Переходим к следующему состоянию
                end
                1: begin 
                    led <= 4'b0010;  // Включаем второй светодиод
                    i <= i + 1;      // Переходим к следующему состоянию
                end
                2: begin 
                    led <= 4'b0100;  // Включаем третий светодиод
                    i <= i + 1;      // Переходим к следующему состоянию
                end
                3: begin 
                    led <= 4'b1000;  // Включаем четвертый светодиод
                    i <= 0;          // Возвращаемся к первому состоянию, чтобы цикл повторился
                end
            endcase
        end
    end

endmodule

/*
 * Пояснения:
 * 1. Сигналы и переменные:
 *    - `nrst`: активный низкий сброс, используется для сброса состояния модуля и сброса всех регистров.
 *    - `clk`: основной тактовый сигнал, который используется для обновления состояния системы.
 *    - `led`: 4-битный выходной сигнал для управления 4 светодиодами.
 *    - `counter`: 32-битный счетчик для деления частоты тактового сигнала `clk`.
 *    - `clk2`: разделенный тактовый сигнал, частота которого ниже, чем у основного сигнала `clk`.
 *    - `i`: 8-битный счетчик для индекса текущего состояния последовательности светодиодов.
 *
 * 2. Делитель тактовой частоты:
 *    - С помощью счетчика `counter` генерируется сигнал `clk2` с более низкой частотой.
 *    - Сигнал `clk2` используется для управления обновлением состояния светодиодов.
 *    - Когда счетчик достигает 1250000, сигнал `clk2` переключается, обеспечивая низкочастотный сигнал для управления светодиодами.
 *
 * 3. Управление светодиодами:
 *    - Светодиоды переключаются поочередно. Каждый новый светодиод включается через один цикл `clk2`.
 *    - Когда значение счетчика `i` достигает 3, оно сбрасывается, и цикл повторяется.
 *
 * 4. Принцип работы:
 *    - Когда модуль сбрасывается (`nrst` = 0), все регистры (включая светодиоды) сбрасываются в нулевое состояние.
 *    - После сброса светодиоды начинают поочередно включаться и выключаться с использованием делителя тактовой частоты.
 *
 * Пояснения используемых конструкций Verilog:
 *
 * 1. `module` и `endmodule`:
 *    - `module` и `endmodule` определяют начало и конец модуля в Verilog. Вся логика дизайна находится между этими ключевыми словами.
 *
 * 2. `input`, `output` и `reg`:
 *    - `input` определяет входные сигналы в модуле. В данном случае, это `nrst` и `clk`.
 *    - `output reg` определяет выходной сигнал, который является регистром (регистры могут хранить данные и быть изменены внутри `always` блоков).
 *    - `reg` указывает, что переменная является регистром, который может хранить состояние между тактами.
 *
 * 3. `always`:
 *    - Блок `always` в Verilog используется для описания поведения, которое должно быть выполнено на каждом такте или в ответ на изменение сигналов.
 *    - В данном коде есть два блока `always`: один для делителя тактовой частоты (`clk2`), а второй для управления светодиодами.
 *    - `@(posedge clk or negedge nrst)` означает, что блок выполняется при каждом положительном фронте сигнала `clk` или при нисходящем фронте сигнала `nrst` (сигнал сброса).
 *    - Важно использовать `posedge` (положительный фронт) или `negedge` (негативный фронт) для синхронизации на тактовых сигналах.
 *
 * 4. Операторы `if`, `else`:
 *    - Оператор `if` используется для выполнения действия, если условие истинно. В данном случае, он проверяет сигнал сброса `nrst` или значение счетчика.
 *    - Оператор `else` выполняет альтернативное действие, если условие не выполняется.
 *
 * 5. Оператор `case`:
 *    - Оператор `case` используется для выбора одного из нескольких возможных состояний на основе значения переменной. В данном случае, `i` используется для определения состояния светодиодов.
 *    - Каждое состояние `i` соответствует включению одного из четырех светодиодов.
 *
 * 6. Оператор присваивания `<=` (non-blocking assignment):
 *    - Внутри блоков `always` мы используем оператор `<=`, чтобы присвоить значения переменным. Это называется "неблокирующим присваиванием" и гарантирует, что значения регистров будут обновляться на следующем такте.
 *    - Это важно, чтобы избежать неправильного порядка обновления значений внутри последовательных операций.
 *
 * 7. Сигналы активного низкого сброса (`nrst`):
 *    - Сигнал сброса используется для инициализации состояния системы. В данном случае, когда сигнал `nrst` активен (низкий), все регистры сбрасываются в ноль, и система возвращается в начальное состояние.
 */

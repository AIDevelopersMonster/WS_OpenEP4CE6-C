// ----------------------------------------------------------------------
// Module     : 8 Push Buttons
// Project    : 8 Push Buttons Demo
// Description: Этот модуль управляет светодиодами на основе состояния кнопок.
//              Используется 8 кнопок (key) и 4 светодиода (led).
//              Каждое нажатие кнопки изменяет состояние светодиодов.
//              Система работает с тактовым сигналом (clk) и асинхронным сбросом (reset).
//              Применяется двоичное представление состояний кнопок для управления светодиодами.
// ----------------------------------------------------------------------
//  GitHub Repository: https://github.com/AIDevelopersMonster/WS_OpenEP4CE6-C/
//  YouTube Playlist: https://www.youtube.com/playlist?list=PLVoFIRfTAAI7-d_Yk6bNVnj4atUdMxvT5
// ------------------------------------------------------------


// Входные и выходные сигналы модуля:
module joystick(
    input clk,            // Тактовый сигнал
    input reset,          // Сигнал сброса
    input [7:0] key,      // 8 кнопок (key), каждая из которых управляет состоянием светодиодов
    output [3:0] led      // 4 светодиода (led), которые изменяются в зависимости от нажатых кнопок
);

// Регистры для управления состоянием светодиодов и счетчика:
reg [3:0] led_reg;      // Регистр для хранения состояния светодиодов
reg [10:0] Count1;      // Счётчик для создания задержки
reg Count;              // Флаг для смены состояния светодиодов с задержкой

// Процесс счёта и смены состояния счетчика:
always @(posedge clk or negedge reset) begin
    if (!reset)               // При сбросе счетчик обнуляется
        Count1 <= 11'd0;
    else if (Count1 == 11'd1999)  // Когда счетчик достигает 1999, меняем состояние флага
        Count = ~Count;
    else
        Count1 <= Count1 + 1'b1; // Иначе увеличиваем счетчик
end

// Процесс управления светодиодами на основе нажатых кнопок:
always @(posedge Count or negedge reset) begin
    if (!reset)                          // При сбросе включаются все светодиоды
        led_reg <= 4'b1111;                // Все светодиоды включены
    else if (key == 8'b11111111_11111110) // Когда нажата кнопка 1 (key[0] = 0)
        led_reg <= 4'b1110;                // Включаем все кроме первого светодиода
    else if (key == 8'b11111111_11111101) // Когда нажата кнопка 2 (key[1] = 0)
        led_reg <= 4'b1101;                // Включаем все кроме второго светодиода
    else if (key == 8'b11111111_11111011) // Когда нажата кнопка 3 (key[2] = 0)
        led_reg <= 4'b1100;                // Включаем все кроме третьего светодиода
    else if (key == 8'b11111111_11110111) // Когда нажата кнопка 4 (key[3] = 0)
        led_reg <= 4'b1011;                // Включаем все кроме четвёртого светодиода
    else if (key == 8'b11111111_11101111) // Когда нажата кнопка 5 (key[4] = 0)
        led_reg <= 4'b1010;                // Включаем все кроме пятого светодиода
    else if (key == 8'b11111111_11011111) // Когда нажата кнопка 6 (key[5] = 0)
        led_reg <= 4'b1001;                // Включаем все кроме шестого светодиода
    else if (key == 8'b11111111_10111111) // Когда нажата кнопка 7 (key[6] = 0)
        led_reg <= 4'b1000;                // Включаем все кроме седьмого светодиода
    else if (key == 8'b11111111_01111111) // Когда нажата кнопка 8 (key[7] = 0)
        led_reg <= 4'b0111;                // Включаем все кроме восьмого светодиода
    else
        led_reg <= led_reg;                // Если не нажата ни одна кнопка, сохраняем текущее состояние
end

// Вывод состояния светодиодов:
assign led = led_reg;

endmodule

// Пояснения:
// - Вход "key" представляет собой 8-битное значение, где каждый бит соответствует одной кнопке.
// - Если кнопка нажата (соответствующий бит равен 0), то меняется состояние светодиодов.
// - Для реализации работы используется двоичная система. Например:
//   key == 8'b11111111_11111110 означает, что только первая кнопка нажата (key[0] = 0), остальные 7 кнопок не нажаты (1).
// - Модуль генерирует сигнал для включения/выключения светодиодов в зависимости от нажатых кнопок.
// - Сигнал "reset" выполняет сброс, возвращая все светодиоды в исходное состояние.
